`include "design.sv"
`include "env_config.svh"
`include "dut_interface.sv"
`include "trans1.svh"
`include "tr_sequence.svh"
`include "tb_sequencer.svh"
`include "tb_driver.svh"
`include "tb_monitor.svh"
`include "tb_scoreboard.svh"
`include "tb_agent.svh"
`include "tb_environment.svh"
`include "base_test.svh"
`include "test.sv"
/*`include "sanity_test.svh"
`include "walk_0_test.svh"
`include "walk_1_test.svh"
`include "full_mem_test.svh"
`include "psel_setup_voil_test.svh"
`include "psel_access_voil_test.svh"
`include "penable_setup_voil_test.svh"
`include "penable_access_voil_test.svh"
`include "pwrite_voil_test.svh"
`include "pwdata_voil_test.svh"
`include "paddr_voil_test.svh"
`include "random_test.svh"
`include "rw_with_idle_test.svh"*/
