class transaction;
        logic PENABLE;
        logic PWRITE;
        logic PSEL;
    rand logic [`ADDRWIDTH-1:0] PADDR;
    rand logic [`DATAWIDTH-1:0] PWDATA;
        logic [`DATAWIDTH-1:0] PRDATA;
        logic PREADY;
	


endclass
